module controlUnit();

endmodule
